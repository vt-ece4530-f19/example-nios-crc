
module platformnioscrc (
	clk_clk,
	hex_export,
	reset_reset_n);	

	input		clk_clk;
	output	[23:0]	hex_export;
	input		reset_reset_n;
endmodule
